** Profile: "SCHEMATIC1-simualareac"  [ c:\users\rares\appdata\roaming\spb_data\cdssetup\workspace\projects\proiectcad\proiectcad-pspicefiles\schematic1\simualareac.sim ] 

** Creating circuit file "simualareac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\rares\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 10MEg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
